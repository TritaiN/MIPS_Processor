`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/16/2020 03:11:42 PM
// Design Name: 
// Module Name: instruction_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instruction_mem(
    input [9:0] read_addr,
    output [31:0] data
    );
    
    reg [31:0] rom [255:0];  
    
    initial  
    begin  
		                                                // instruction           alu result            register content       mem content
														
        rom[0] = 32'b00100000001000010000000000000110; // addi r1,r0,#6             6; b110; d6                r1=6                   -
//        rom[1] = 32'b11000000001000000000100010000000; // sll r1, r1, 2             b11000, d24                 r1 = 24         
//        rom[2] = 32'b00110000001000100000000000000000; //andi r1, r2, 2             b0, d0                 r2 = d0
//        rom[3] = 32'b00000000010000010000000000100111;  //nor r2, r1, r0             b00100, d8                  r0 = 8 
//        rom[4] = 32'b00000000000000010000100000101010; //slt r0, r1, r1             b1, d1                      r1 = 1
//        rom[5] = 32'b00100000010000100000000000000111; //addi r2, r2, 3             d3                          r2 = 7
//        rom[6] = 32'b11000000010000000001100010000010; //srl r2, r3, 2            b1, d1                       r3 = 1 
//        rom[7] = 32'b11000000001000010000111111000000; // sll r1, r1, 31             b111..00,                 r1 = 11..00
//        rom[8] = 32'b11000000001000000000001111000011; //sra r1, r1,31             b01                         r1 = 1
//        rom[9] = 32'b00000000011000100001000000100110; //xor r3, r2, r2            d6, b001100                  r2 = d6
//        rom[10]=  32'b00100000100001000000000000000010; // addi r4,r4,#2             2; b10; d2                r4=2        
//        rom[11] = 32'b00000000010001000010100000011000;//mult r2, r4, r4                                      
//        rom[12] = 32'b00000000010001010001100000011010; //div r2, r3, r2            
//        rom[13] = 32'b00010000001000000000000000000010; //beq 
//        rom[14] = 32'b00010000110001110000000000000001; //beq 
//        rom[15] = 32'b11000000001000000000001111000011; // skipping because of branch
//        rom[16] = 32'b00001000000000000000000000010011; //jump to instruction 19
//        rom[17] = 32'b00100000000000010000000000000111; //   
//        rom[18] = 32'b11000000001000000000100010000000; //   
//        rom[19] = 32'b00100000000000010000000000001111; // addi r1,r0,#15             15; b1111;                 r1=15     
        //rom[20] = 32'b00100000000000010000000000011111; // addi r1,r0,#31             15; b11111;                 r1=31   
        /*rom[1]  = 32'b00100000000000100000000000001110; // addi r2,r0,#e                 e                    r2=e                   -
        rom[2]  = 32'b00100000000000110000000001001110; // addi r3,r0,#4e                4e                   r3=4e                  -
        rom[3]  = 32'b00100000000001000000000011010010; // addi r4,r0,#d2                d2                   r4=d2                  -
        rom[4]  = 32'b00100000000001011110000110010101; // addi r5,r0,#e195           ffffe195                r5=ffffe195            -
        rom[5]  = 32'b00100000000001101111111000010010; // addi r6,r0,#fe12           fffffe12                r6=fffffe12            -
        rom[6]  = 32'b00000000001001000011100000100000; // add r7,r1,r4                  d8                   r7=d8                  -
        rom[7]  = 32'b00000000011001010100000000100000; // add r8,r3,r5               ffffe1e3                r8=ffffe1e3            -
        rom[8]  = 32'b10101100001001110000000000000010; // sw mem[r1+2] <= r7            8                    -                   mem[2]=d8
        rom[9]  = 32'b10101100100010001111111111111110; // sw mem[r4-2] <= r8            d0                   -                   mem[52]=ffffe1e3
        rom[10] = 32'b00000000100000100100100000100010; // sub r9,r4,r2                  C4                   r9=c4                  -
        rom[11] = 32'b00000000001001010101000000100010; // sub r10,r1,r5                1e71                  r10=1e71               -
        rom[12] = 32'b10101101001010100000000000000000; // sw mem[r9+0] <= r10           c4                   -                   mem[49]=1e71
        rom[13] = 32'b00000001001001110101100000100101; // or r11,r9,r7                  dc                   r11=dc                 -
        rom[14] = 32'b00000001000010100110000000100100; // and r12,r8,r10                61                   r12=61                 -
        rom[15] = 32'b10001100001011010000000000000010; // r13 =mem[r1+2]                8                    r13=d8                 -
        rom[16] = 32'b10001100100011101111111111111110; // r14 =mem[r4-2]                d0                   r14=ffffe1e3           -
        rom[17] = 32'b10001101001011110000000000000000; // r15 =mem[r9+0]                c4                   r15=1e71               - 
        */   
      end  
      
      assign data = rom[read_addr[9:2]];

endmodule
